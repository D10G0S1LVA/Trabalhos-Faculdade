* C:\Users\Diogo Silva\Desktop\VideoEscola\EA\Lab1_exerc6.sch

* Schematics Version 9.1 - Web Update 1
* Wed Apr 15 20:50:55 2020



** Analysis setup **
.tran 0ns 60ms 0 10000ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Lab1_exerc6.net"
.INC "Lab1_exerc6.als"


.probe


.END
