* D:\VideoEscola\Eletronica Analogica\Lab4 transistores.sch

* Schematics Version 9.2
* Thu Jun 04 16:12:41 2020



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Lab4 transistores.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
