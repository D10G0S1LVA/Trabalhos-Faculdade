* D:\VideoEscola\Eletronica Analogica\Lab5 3 exercicio1.sch

* Schematics Version 9.2
* Tue Jul 07 15:33:33 2020



** Analysis setup **
.OP 
.LIB "D:\VideoEscola\Eletronica Analogica\Lab5 3 exercicio1.lib"


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Lab5 3 exercicio1.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
