* D:\VideoEscola\Eletronica Analogica\Lab5 2 exercicio.sch

* Schematics Version 9.2
* Tue Jul 07 18:47:35 2020



** Analysis setup **
.OP 
.LIB "D:\VideoEscola\Eletronica Analogica\Lab5 2 exercicio.lib"


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Lab5 2 exercicio.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
