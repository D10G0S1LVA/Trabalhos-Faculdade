* C:\Users\joaoq\Desktop\lixo\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Tue Jun 16 16:49:08 2020



** Analysis setup **
.DC LIN V_VCC 0 +10 0.01 
+ OCT V_VBB 2.7 10.7 2 
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
