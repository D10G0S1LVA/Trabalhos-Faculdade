* D:\VideoEscola\Eletronica Analogica\Lab5 4 exercicio1.sch

* Schematics Version 9.2
* Mon Jul 06 15:41:26 2020



** Analysis setup **
.OP 
.LIB "D:\VideoEscola\Eletronica Analogica\Lab5 4 exercicio1.lib"


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Lab5 4 exercicio1.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
