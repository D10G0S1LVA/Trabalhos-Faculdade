* D:\VideoEscola\Eletronica Analogica\Lab5 4 exercicio.sch

* Schematics Version 9.2
* Mon Jul 06 14:48:54 2020



** Analysis setup **
.OP 
.LIB "D:\VideoEscola\Eletronica Analogica\Lab5 4 exercicio.lib"


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Lab5 4 exercicio.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
