* D:\VideoEscola\Eletronica Analogica\Lab5 3 exercicio.sch

* Schematics Version 9.2
* Mon Jul 06 13:16:37 2020



** Analysis setup **
.OP 
.LIB "D:\VideoEscola\Eletronica Analogica\Lab5 3 exercicio.lib"


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Lab5 3 exercicio.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
