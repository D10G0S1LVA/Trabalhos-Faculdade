* D:\VideoEscola\Eletronica Analogica\Lab5 5 exercicio.sch

* Schematics Version 9.2
* Tue Jul 07 20:48:07 2020



** Analysis setup **
.tran 0ns 2.6
.OP 
.LIB "D:\VideoEscola\Eletronica Analogica\Lab5 5 exercicio.lib"


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Lab5 5 exercicio.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
