* C:\Users\Diogo Silva\Desktop\VideoEscola\EA\Lab1_exerc8.sch

* Schematics Version 9.1 - Web Update 1
* Wed Apr 15 20:41:54 2020



** Analysis setup **
.tran 0ns 20s 0 1000ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Lab1_exerc8.net"
.INC "Lab1_exerc8.als"


.probe


.END
